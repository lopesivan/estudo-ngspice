# exemplo de operação com let

.control
let myvector = [1, 2, 3, 4, 5]
let newvector = myvector + 1
.endc

.end

