.param Vvalue  = 25V           ; tensão fornecida
.param Rvalue  = 1.2Meg        ; valor da resistência
.param Cvalue  = 20uF          ; valor da Capacitância
.param tau     = Rvalue*Cvalue

** circuito:
*         1         2
* v_i(t) ---[ R ]---+---[ C ]--- GND
*                   |
*               v_out(t)
*

V0 n1 GND  PULSE(0 {Vvalue} 1u 1u 1u 1   1)
* V0 n1 GND  PULSE(0 {Vvalue} 0  1u 1u 1m 2m)
R1 n1  n2  {Rvalue}
C1 n2 GND  {Cvalue}
