.tran {tau/1000} {5*tau}
