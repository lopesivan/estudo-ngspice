Exemplo de operações com Complexos

.control
    let z1 = (4, 5)
    let z2 = (1, -2)
    print z1
    print z2
    let r = z1+z2
    print r
    print real(r)
    print imag(r)
    print phase(r)
    set units = degrees
    print phase(r)
.endc

.end
